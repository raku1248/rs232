
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Receiver is
end Receiver;

architecture Behavioral of Receiver is

begin


end Behavioral;

